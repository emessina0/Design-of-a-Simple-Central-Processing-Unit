library verilog;
use verilog.vl_types.all;
entity Processor3_vlg_vec_tst is
end Processor3_vlg_vec_tst;
