library verilog;
use verilog.vl_types.all;
entity Processor2_vlg_vec_tst is
end Processor2_vlg_vec_tst;
